package classes_pkg;
  `include "Transaction.sv"
  `include "Generator.sv"
  `include "Driver.sv"
  `include "Monitor.sv"
  `include "Scoreboard.sv"
  `include "Environment.sv"
  
endpackage
